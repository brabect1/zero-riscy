package zeroriscy_pkg;

    typedef logic[33:0] t_instr;

    localparam int irq = 32;
    localparam int dirq = 33;

endpackage: zeroriscy_pkg
